module main

// import year_2023.day_1.part_1
// import year_2023.day_1.part_2
// import year_2023.day_2.part_1
import year_2023.day_2

fn main() {
	// println(part_1.solve(part_1.actual_input))
	// println(part_2.solve(part_2.actual_input))
	// assert part_1.solve(part_1.example_input) == part_1.example_output
	assert day_2.part_1(day_2.example_input) == day_2.example_output_part_1
	println(day_2.part_1(day_2.input))
	assert day_2.part_2(day_2.example_input) == day_2.example_output_part_2
	println(day_2.part_2(day_2.input))
}
