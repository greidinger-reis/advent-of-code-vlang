module main

// import year_2023.day_1.part_1
import year_2023.day_1.part_2

fn main() {
	dump(part_2.solve(part_2.actual_input))
}
