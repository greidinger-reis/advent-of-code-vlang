module main

// import year_2023.day_1.part_1
// import year_2023.day_1.part_2
import year_2023.day_2.part_1

fn main() {
	// println(part_1.solve(part_1.actual_input))
	// println(part_2.solve(part_2.actual_input))
    part_1.solve(part_1.example_input)
}
