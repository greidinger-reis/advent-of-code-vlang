module main

import day_3

fn main() {
	println(day_3.part_2(day_3.input))
}
