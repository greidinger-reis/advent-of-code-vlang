module main

import day_4

fn main() {
	println(day_4.part_2(day_4.input))
}
