module main

import day_5

fn main() {
	println(day_5.part_1(day_5.input))
}
